noise_1
V1 N005 0 V value=0 dc=0 dcvar=0 noise=0
R1 N001 N005 R value={R_s} noisetemp={T} noiseflow=0 dcvar=0 dcvarlot=0
I1 N004 0 I value=0 dc=0 dcvar=0 noise={4*k*T*n*Gamma*g_m}
H1 N003 in N004 N006 {1/g_m}
F1 in 0 N006 0 {s/(2*pi*f_T)}
V2 N003 N002 V value=0 dc=0 dcvar=0 noise={4*k*T*n*Gamma*f_ell^AF/g_m/f}
L1 N001 N002 L value={L_s} iinit=0
E1 out 0 in 0 {1/(s*tau_i)}
R2 N002 0 R value={R_t} noisetemp={T} noiseflow=0 dcvar=0 dcvarlot=0
.param f_ell={alpha*f_T^(1/AF)} f_T={g_m/(2*pi*c_iss)}
.param n=1.35 Gamma={2/3} AF=1 alpha=0.0033
.param L_s = 120m R_s=875 tau_i=15.9u
.param R_t=10k
* Rceive coil (resonance  not modeled > 150 kHz)
* Shot noise associated with the DC gate current is not modeled (IG = 0)
* Channel current noise
* Input-referred flicker noise
* Gate-\ninduced\nnoise
* Input-\nreferred\nchannel\nvoltage\nnoise
* Integrating voltage amplifier
* Termination resistor
.end
